// ********************************************************************
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// ********************************************************************
// File name    : clk_tb.v
// Module name  : clk_tb
// Author       : 薛骏
// Description  : 用于仿真时钟分频模块波形
// 
// --------------------------------------------------------------------
// Code Revision History : 
// --------------------------------------------------------------------
// Version: |Mod. Date:
// V1.0     |2019/12/10
// --------------------------------------------------------------------
// Module Function: 模块波形仿真

`timescale 1ns / 100ps
module clk_tb;

	reg clki;
	wire clk_out;
	
	// 设置时钟信号
	parameter CLOCK = 20;
	initial
		clki = 0;
	always
		#(CLOCK) clki = ~clki;
	
	// 例化模块（以5分频为例）
	clk #(.num(10_000_000)) c1(.clk(clki),
			 .clkout(clk_out));

endmodule
